`timescale 1ns / 1ps


module Mealy1101(clk, rst, data, out);

    input clk, rst, data;
    output out;
    reg [3:0] temp;
    reg out;
    
    
    initial temp = 4'b0000;
    initial out = 1'b0;
        
        always @(posedge clk)begin
        temp =(temp << 1)+data;
        
        if(rst == 1'b1) begin
        temp = 4'b0000;
        out = 1'b0;
        end
        
        else if(temp ==4'b1101) out =1'b1;
        else out = 1'b0;
        
        end
    
endmodule
