`timescale 1ns / 1ps


module conver(
    input a, b, c, d,
    output e, f, g, h
    );
    
    assign e = ~(~(a&a)&~(~(~(~(~(b&d)&~(b&d))&~(~(b&d)&~(b&d)))&~(~(~(b&c)&~(b&c))&~(~(b&c)&~(b&c))))&~(~(~(~(b&d)&~(b&d))&~(~(b&d)&~(b&d)))&~(~(~(b&c)&~(b&c))&~(~(b&c)&~(b&c))))));
    assign f = ~(~(a&a)&~(~(~(~(~(b&c)&~(b&c))&~(~(b&c)&~(b&c)))&~(~(~(b&~d)&~(b&~d))&~(~(b&~d)&~(b&~d))))&~(~(~(~(b&c)&~(b&c))&~(~(b&c)&~(b&c)))&~(~(~(b&~d)&~(b&~d))&~(~(b&~d)&~(b&~d))))));
    assign g = ~(~(a&a)&~(~(~(~(~(~(~(b&~c)&~(b&~c))&d)&~(~(~(b&~c)&~(b&~c))&d))&~(~(~(~(b&~c)&~(b&~c))&d)&~(~(~(b&~c)&~(b&~c))&d)))&~(~(~(~b&c)&~(~b&c))&~(~(~b&c)&~(~b&c))))&~(~(~(~(~(~(b&~c)&~(b&~c))&d)&~(~(~(b&~c)&~(b&~c))&d))&~(~(~(~(b&~c)&~(b&~c))&d)&~(~(~(b&~c)&~(b&~c))&d)))&~(~(~(~b&c)&~(~b&c))&~(~(~b&c)&~(~b&c))))));
    assign h = d;

    
endmodule
